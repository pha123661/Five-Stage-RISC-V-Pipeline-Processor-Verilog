module Hazard_detection(
input [4:0] IFID_regRs,
input [4:0] IFID_regRt,
input [4:0] IDEXE_regRd,
input IDEXE_memRead,
output PC_write,
output IFID_write,
output control_output_select
);


endmodule

